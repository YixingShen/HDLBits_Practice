module top_module (
    input [7:0] a, b, c, d,
    output [7:0] min);//

    // assign intermediate_result1 = compare? true: false;
    
    always @(*) begin
        min = a;

        if (b < min) min = b;
        if (c < min) min = c;
        if (d < min) min = d;
    end

endmodule