//The following adder-subtractor with zero flag doesn't work. Fix the bug(s).

//// synthesis verilog_input_version verilog_2001
//module top_module ( 
//    input do_sub,
//    input [7:0] a,
//    input [7:0] b,
//    output reg [7:0] out,
//    output reg result_is_zero
//);//
//
//    always @(*) begin
//        case (do_sub)
//          0: out = a+b;
//          1: out = a-b;
//        endcase
//
//        if (~out)
//            result_is_zero = 1;
//    end
//
//endmodule

// synthesis verilog_input_version verilog_2001
module top_module ( 
    input do_sub,
    input [7:0] a,
    input [7:0] b,
    output reg [7:0] out,
    output reg result_is_zero
);//

    always @(*) begin
        case (do_sub)
          0: out = a+b;
          1: out = a-b;
        endcase

        result_is_zero = (out == 0) ? 1 : 0;
 
    end

endmodule