module top_module (
    input clk,
    input d, 
    input ar,   // asynchronous reset
    output reg q);

    always @(posedge clk, posedge ar) begin
        if (ar == 1) begin
            q <= 0;
        end
        else begin
            q <= d;
        end
    end

endmodule
