//You are provided with a BCD one-digit adder named bcd_fadd that adds two BCD digits and carry-in, and produces a sum and carry-out.
//
//module bcd_fadd {
//    input [3:0] a,
//    input [3:0] b,
//    input     cin,
//    output   cout,
//    output [3:0] sum );
//Instantiate 100 copies of bcd_fadd to create a 100-digit BCD ripple-carry adder. Your adder should add two 100-digit BCD numbers
// (packed into 400-bit vectors) and a carry-in to produce a 100-digit sum and carry out.

//Hint...
//An instance array or generate statement would be useful here.

module top_module( 
    input [399:0] a, b,
    input cin,
    output cout,
    output [399:0] sum );

    wire [99:0] cout_t;

    bcd_fadd inst(.a(a[3:0]),
              .b(b[3:0]),
              .cin(cin),
              .cout(cout_t[0]),
              .sum(sum[3:0]));
              
    genvar i;
    generate
        for (i = 1; i < 100; i++) begin: myForLoop
            bcd_fadd inst(.a(a[3+i*4:i*4]),
                          .b(b[3+i*4:i*4]),
                          .cin(cout_t[i - 1]),
                          .cout(cout_t[i]),
                          .sum(sum[3+i*4:i*4]));
        end
    endgenerate

    assign cout = cout_t[99];
    
endmodule
